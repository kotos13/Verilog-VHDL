/*--------------------------------------------------------------------------------
Module Name:    CPLD_CONTROL_tb_func
--------------------------------------------------------------------------------*/

`timescale	1 ps / 1 ps

module CPLD_CONTROL_tb_func

endmodule
